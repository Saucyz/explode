-- Inputs: SW7°0 are parallel port inputs to the Nios II system.
-- CLOCK_50 is the system clock.
-- KEY0 is the active-low system reset.
-- Outputs: LEDG7°0 are parallel port outputs from the Nios II system.
-- SDRAM ports correspond to the signals in Figure 2; their names are those
-- used in the DE2 User Manual.
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;
USE ieee.std_logic_unsigned.all;

ENTITY Mod2 IS

PORT (
	SW : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	KEY : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	CLOCK_50 : IN STD_LOGIC;
	
	LEDG : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);

	UART_RXD           : in    std_logic;             -- RXD
   UART_TXD           : out   std_logic;             -- TXD

	DRAM_CLK, DRAM_CKE : OUT STD_LOGIC;
	DRAM_ADDR : OUT STD_LOGIC_VECTOR(11 DOWNTO 0);
	DRAM_BA_0, DRAM_BA_1 : BUFFER STD_LOGIC;
	DRAM_CS_N, DRAM_CAS_N, DRAM_RAS_N, DRAM_WE_N : OUT STD_LOGIC;
	DRAM_DQ : INOUT STD_LOGIC_VECTOR(15 DOWNTO 0);
	DRAM_UDQM, DRAM_LDQM : BUFFER STD_LOGIC;

	LCD_DATA : inout STD_LOGIC_VECTOR(7 downto 0);
	LCD_ON, LCD_BLON, LCD_EN, LCD_RS, LCD_RW : out STD_LOGIC;
	
	SD_CMD, SD_DAT, SD_DAT3 : INOUT STD_LOGIC;
	SD_CLK : OUT STD_LOGIC;
	
	AUD_ADCDAT         : in    std_logic;             -- ADCDAT
	AUD_ADCLRCK        : in    std_logic;             -- ADCLRCK
   AUD_BCLK           : in    std_logic;             -- BCLK
   AUD_DACDAT         : out   std_logic;             -- DACDAT
   AUD_DACLRCK        : in    std_logic;             -- DACLRCK
	
	I2C_SDAT    : inout std_logic;
	I2C_SCLK    : out   std_logic;
	
	CLOCK_27	:	IN STD_LOGIC;
	AUD_XCK	:	OUT STD_LOGIC;
	TD_RESET : OUT STD_LOGIC
	);
	
END Mod2;

ARCHITECTURE Structure OF Mod2 IS
COMPONENT nios_system
PORT (
	clk_clk : IN STD_LOGIC;
	reset_reset_n : IN STD_LOGIC;
	
	sdram_clk_clk : OUT STD_LOGIC;
	
	leds_export : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
	switches_export : IN STD_LOGIC_VECTOR(7 DOWNTO 0);

	serial_RXD           : in    std_logic                     := 'X';             -- RXD
   serial_TXD           : out   std_logic;                                        -- TXD
	
	sdram_wire_addr : OUT STD_LOGIC_VECTOR(11 DOWNTO 0);
	sdram_wire_ba : BUFFER STD_LOGIC_VECTOR(1 DOWNTO 0);
	sdram_wire_cas_n : OUT STD_LOGIC;
	sdram_wire_cke : OUT STD_LOGIC;
	sdram_wire_cs_n : OUT STD_LOGIC;
	sdram_wire_dq : INOUT STD_LOGIC_VECTOR(15 DOWNTO 0);
	sdram_wire_dqm : BUFFER STD_LOGIC_VECTOR(1 DOWNTO 0);
	sdram_wire_ras_n : OUT STD_LOGIC;
	sdram_wire_we_n : OUT STD_LOGIC;
	
	lcd_data_DATA : INOUT STD_LOGIC_VECTOR(7 downto 0);
	lcd_data_ON : OUT STD_LOGIC;
	lcd_data_BLON : OUT STD_LOGIC;
	lcd_data_EN : OUT STD_LOGIC;
	lcd_data_RS : OUT STD_LOGIC;
	lcd_data_RW : OUT STD_LOGIC;
	
	keys_export : IN STD_LOGIC_VECTOR(3 downto 0);
	
	sd_wire_b_SD_cmd   : inout std_logic := 'X';             -- b_SD_cmd
   sd_wire_b_SD_dat   : inout std_logic := 'X';             -- b_SD_dat
   sd_wire_b_SD_dat3  : inout std_logic := 'X';             -- b_SD_dat3
   sd_wire_o_SD_clock : out   std_logic;                     -- o_SD_clock
		
	audio_ADCDAT         : in    std_logic                     := 'X';             -- ADCDAT
	audio_ADCLRCK        : in    std_logic                     := 'X';             -- ADCLRCK
   audio_BCLK           : in    std_logic                     := 'X';             -- BCLK
   audio_DACDAT         : out   std_logic;                                        -- DACDAT
   audio_DACLRCK        : in    std_logic                     := 'X';             -- DACLRCK
	
	audio_config_SDAT    : inout std_logic                     := 'X';             -- SDAT
   audio_config_SCLK    : out   std_logic;                                        -- SCLK
	
	audio_clk_clk				:	OUT STD_LOGIC;
	clk_in_secondary_clk		:	IN STD_LOGIC
	);
END COMPONENT;

SIGNAL DQM : STD_LOGIC_VECTOR(1 DOWNTO 0);
SIGNAL BA : STD_LOGIC_VECTOR(1 DOWNTO 0);

BEGIN
DRAM_BA_0 <= BA(0);
DRAM_BA_1 <= BA(1);
DRAM_UDQM <= DQM(1);
DRAM_LDQM <= DQM(0);
 TD_RESET <= '1';

-- Instantiate the Nios II system entity generated by the Qsys tool.
NiosII: nios_system
PORT MAP (
	clk_clk => CLOCK_50,
	reset_reset_n => KEY(0),
	
	sdram_clk_clk => DRAM_CLK,
	
	leds_export => LEDG,
	switches_export => SW,
	
	serial_RXD => UART_RXD,
	serial_TXD => UART_TXD,

	sdram_wire_addr => DRAM_ADDR,
	sdram_wire_ba => BA,
	sdram_wire_cas_n => DRAM_CAS_N,
	sdram_wire_cke => DRAM_CKE,
	sdram_wire_cs_n => DRAM_CS_N,
	sdram_wire_dq => DRAM_DQ,
	sdram_wire_dqm => DQM,
	sdram_wire_ras_n => DRAM_RAS_N,
	sdram_wire_we_n => DRAM_WE_N,

	lcd_data_DATA => LCD_DATA,
	lcd_data_ON => LCD_ON,
	lcd_data_BLON => LCD_BLON,
	lcd_data_EN => LCD_EN,
	lcd_data_RS => LCD_RS,
	lcd_data_RW => LCD_RW,
	
	keys_export => KEY,
	
	sd_wire_b_SD_cmd   => SD_CMD,   --    			sd_wire.b_SD_cmd
   sd_wire_b_SD_dat   => SD_DAT,   --           .b_SD_dat
   sd_wire_b_SD_dat3  => SD_DAT3,  --           .b_SD_dat3
   sd_wire_o_SD_clock => SD_CLK,   --           .o_SD_clock
		
	audio_ADCDAT 			=> AUD_ADCDAT,
	audio_ADCLRCK 			=> AUD_ADCLRCK,
	audio_BCLK    			=> AUD_BCLK,
	audio_DACDAT  			=> AUD_DACDAT,
	audio_DACLRCK 			=> AUD_DACLRCK,
	
	audio_config_SDAT    => I2C_SDAT,    --   audio_config.SDAT
   audio_config_SCLK    => I2C_SCLK,    --               .SCLK
	
	clk_in_secondary_clk	=>	CLOCK_27,
	audio_clk_clk	=>	AUD_XCK
	);

	--DRAM_CLK <= CLOCK_50;
END Structure;